module CP
(
input clk, in, rst, in_sop,
input signed [19:0] in_i, in_q,
output out_sop,
output signed [19:0] out_i, out_q
);









endmodule
